module FloatingPointAddition();

input logic [31:0] a;
input logic [31:0] b;
input logic start;
output logic [31:0] result;
output logic valid;
output logic ready;



import floatingpoint::*;


	
endmodule